library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
use unisim.vcomponents.all;
--
------------------------------------------------------------------------------------
--
-- Main Entity for ring_osc
--
entity ring_osc is
    port(   Output_clock    : out std_logic;
            previous_sig    : in std_logic;
            ColEN           : in std_logic;
            RowEN           : in std_logic );
end ring_osc;
--
------------------------------------------------------------------------------------
-- 
-- Start of Main Architecture for ring_osc
--	 
architecture low_level_definition of ring_osc is
--
    signal ring_delay1      : std_logic;
    signal ring_delay2      : std_logic;
    signal ring_delay3      : std_logic;
    signal ring_delay4      : std_logic;
    signal ring_invert      : std_logic;
    signal clk_div2         : std_logic;
    signal reset            : std_logic;
    signal toggle           : std_logic;

--
-- Attributes to stop delay logic from being optimised.
--
    attribute dont_touch                : string; 
    attribute dont_touch of ring_delay1 : signal is "true"; 
    attribute dont_touch of ring_delay2 : signal is "true"; 
    attribute dont_touch of ring_delay3 : signal is "true"; 
    attribute dont_touch of ring_delay4 : signal is "true";     
    attribute dont_touch of ring_invert : signal is "true";
    
    attribute dont_touch of Xor_out     : label is "true";
    attribute dont_touch of div2_lut    : label is "true";
    

----all in one slice
    attribute RLOC                  : string;
    attribute RLOC of delay1_lut    : label  is "X0Y0";
    attribute RLOC of delay2_lut    : label  is "X0Y0";
    attribute RLOC of delay3_lut    : label  is "X0Y0";
    attribute RLOC of delay4_lut    : label  is "X0Y0";
    attribute RLOC of div2_lut      : label  is "X0Y0";
    attribute RLOC of En_row_col    : label  is "X0Y0";
    attribute RLOC of invert_lut    : label  is "X0Y0";
    attribute RLOC of Xor_out       : label  is "X0Y0";
    attribute RLOC of toggle_flop   : label  is "X0Y0";

--assign position of all cells
    attribute BEL                   : string;
    attribute BEL of delay1_lut     : label  is "D6LUT";
    attribute BEL of delay2_lut     : label  is "D5LUT";
    attribute BEL of delay3_lut     : label  is "C6LUT";
    attribute BEL of delay4_lut     : label  is "C5LUT";
    attribute BEL of invert_lut     : label  is "B5LUT";
    attribute BEL of Xor_out        : label  is "B6LUT";
    attribute BEL of div2_lut       : label  is "A5LUT";
    attribute BEL of En_row_col     : label  is "A6LUT";
    attribute BEL of toggle_flop    : label  is "BFF";

------------------------------------------------------------------------------------
--	
-- Circuit description
--
------------------------------------------------------------------------------------
--	
begin
--
--Output is the ring oscillator divided by 8 to provide a square wave.
--4 flipflop to divide the signal 8 times

--This LUT is A NAND gate to enable or disable all ring oscillator
En_row_col: component LUT2
    generic map(    INIT    => X"7")
    port map(       I0      => ColEN,
                    I1      => RowEN,
                    O       => reset);
--This LUT is a XOR.  XOR the signal generated by the RO before, 
--in order to receive only one output at the end. 
Xor_out: component LUT2
    generic map(    INIT    => X"6")
    port map(       I0      => clk_div2,
                    I1      => previous_sig,
                    O       => Output_clock);
--to divide the clock   
toggle_flop: component FD
    port map(   D   => toggle,
                Q   => clk_div2,
                C   => ring_invert);

div2_lut: component LUT1
    generic map(    INIT    => X"1")
    port map(       I0      => clk_div2,
                    O       => toggle);
--
--Ring oscillator is formed of 5 delays, all of which are inverters.
-- the other 4 are just used as delay
--
delay1_lut: component LUT1
    generic map(    INIT    => X"1")
    port map(       I0      => ring_invert,
                    O       => ring_delay1);

delay2_lut: component LUT1
    generic map(    INIT    => X"1")
    port map(       I0      => ring_delay1,
                    O       => ring_delay2);

delay3_lut: component LUT1
    generic map(    INIT    => X"1")
    port map(       I0      => ring_delay2,
                    O       => ring_delay3);

delay4_lut: component LUT1
    generic map(    INIT    => X"1")
    port map(       I0      => ring_delay3,
                    O       => ring_delay4 );

invert_lut: component LUT2
    generic map(    INIT    => X"B") 
    port map(       I0      => reset,
                    I1      => ring_delay4,
                    O       => ring_invert );
end low_level_definition;
